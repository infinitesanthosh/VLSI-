Write a Verilog module using a continuous assignment to implement out = a & b.
